-- vhdl-linter-disable type-resolved
LIBRARY IEEE;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY FCS_parallel IS

PORT(
    CLK : IN STD_LOGIC
);

END FCS_parallel;

architecture rtl of  FCS_parallel is

    begin

END architecture rtl;
